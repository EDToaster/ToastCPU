import mem_write_data_source_t::*;
import mem_write_addr_source_t::*;