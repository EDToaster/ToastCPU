
module clock (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
