module datapath (
	
	

);

endmodule